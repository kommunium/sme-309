//`timescale 1ns/1ps
`include "../src/ALU.v"

module ALU_tb();

  reg [31:0] A;
  reg [31:0] B;
  reg [1:0] ALUControl;
  wire [31:0] Result;
  wire [3:0] ALUFlags;

  initial
    begin
      #0 A = 32'b11111111111111111111111111111111;
      B = 32'b11111111111111111111111111111111;
      ALUControl = 2'b00;
      #5 A = 32'b00010000000000000000000000000000;
      B = 32'b00100000000000000000000000000000;
      ALUControl = 2'b00;
      #5 A = 32'b10100000000000000000000000000000;
      B = 32'b10010000000000000000000000000000;
      ALUControl = 2'b00;
      #5 A = 32'b00100000000000000000000000000000;
      B = 32'b01110000000000000000000000000000;
      ALUControl = 2'b00;
      #5 A = 32'b11110000000000000000000000000000;
      B = 32'b00100000000000000000000000000000;
      ALUControl = 2'b00;
      #5 A = 32'b00000000000000000000000000000000;
      B = 32'b00000000000000000000000000000000;
      ALUControl = 2'b00;
      #5 A = 32'b00010000000000000000000000000000;
      B = 32'b11110000000000000000000000000000;
      ALUControl = 2'b00;
      #5 A = 32'b00010000000000000000000000000000;
      B = 32'b00010000000000000000000000000000;
      ALUControl = 2'b01;
      #5 A = 32'b00100000000000000000000000000000;
      B = 32'b00010000000000000000000000000000;
      ALUControl = 2'b01;
      #5 B = 32'b00100000000000000000000000000000;
      A = 32'b00010000000000000000000000000000;
      ALUControl = 2'b01;
    end

  ALU ALU1(
        A,
        B,
        ALUControl,
        Result,
        ALUFlags
      );

endmodule
