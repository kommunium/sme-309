module Multiplier(
    input CLK_MUL, //! dedicated clock signal for multicycle multiply, the frequency is much higher than the CPU clock.
    input Reset, //!  Connect this to the reset of the ARM processor.
    input MUL_EN, //! Multi-cycle Enable. The control unit should assert this when an instruction with a multi-cycle operation is detected
    input MULOp, //! Multi-cycle Operation. "high" for signed multiplication, "low" for unsigned multiplication, Generated by Control unit
    input [31:0] Operand1, //! Multiplicand A
    input [31:0] Operand2, //! Multiplier B

    input [31:0] Sum, //! Provides interface to the 32bit Fulladder in ALU
    output [31:0] MAddInA, //! Provides interface to the 32bit Fulladder in ALU
    output [31:0] MAddInB,
    output MCin, //! Provides interface to the 32bit Fulladder in ALU

    output [31:0] Result, //! LSW(Least Significant Word) of the Product
    output reg Busy //! Set immediately when Start is set. Cleared when the Results become ready. This bit can be used to stall the processor while multi-cycle operations are on.(i.e. keep the PC from fetching next instruction if the multicycle multiply is not finished)
  );

  reg [5:0] counter;
  //! Initialize
  always @(*)
    if(~MUL_EN | Reset)
      begin
        Busy <= 0'b0;
        counter <= 6'b000000;
      end

  reg [63:0] Product;
  //! Detect the start of the multiplication
  always @(posedge CLK_MUL)
    if (MUL_EN & ~Busy & ~counter[5])
      begin
        Busy <= 0'b1;
        Product <= {{32'b0}, Operand2};
        counter <= 6'b000000;
      end


  //! Detect the end of the multiplication
  always @(*)
    if (counter[5])
      Busy <= 0'b0;

  //! Do multiplication
  always @(posedge CLK_MUL)
    if (MUL_EN & Busy)
      begin
        Product <= {{MULOp & Operand1[31]}, Sum, Product[31:1]};
        counter <= counter + 6'b000001;
      end

  //!  Defines the partial product
  assign MAddInA = Product[63:32];
  assign MAddInB = ({32{&counter[4:0] & MULOp & Operand2[31]}}) ^ (Operand1 & {32{Product[0]}});
  assign MCin = &counter[4:0] & MULOp & Operand2[31];
  assign Result = Product[31:0];

endmodule
